.param a=1
.param b=2
.param c=3
.param d=4
.param e=5
.param f=6
