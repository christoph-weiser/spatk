.param a = 1
.param b = 2
.param c = 3
+ d = 4 
+ e = 5
.param f = 6
